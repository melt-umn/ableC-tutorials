grammar edu:umn:cs:melt:tutorials:ableC:intconst:concretesyntax;

imports edu:umn:cs:melt:ableC:concretesyntax;
imports silver:langutil only ast; 

imports edu:umn:cs:melt:tutorials:ableC:intconst:abstractsyntax;

exports edu:umn:cs:melt:tutorials:ableC:intconst:concretesyntax:decl;
exports edu:umn:cs:melt:tutorials:ableC:intconst:concretesyntax:ref;
